3 4
4 1 2 0 3
2 1 3
5 1 3 0 0 2